/cad/dk/PDK_CRN45GS_DGO_11_25/digital/Back_End/lef/tpbn45v_ds_150a/wb/8m/8M_5X2Z/lef/tpbn45v_ds_8lm.lef