/cad/dk/PDK_CRN45GS_DGO_11_25/digital/Back_End/lef/tpfn40lpgv2od3_120a/mt_2/8lm/lef/antenna_8lm.lef