/cad/dk/PDK_CRN45GS_DGO_11_25/IMEC_RAM_generator/ram/ts1n40lpb4096x32m4m_250a/LEF/ts1n40lpb4096x32m4m_250a_4m.lef